module my_module;
endmodule